module controller (
    input clk, rst,
	input[3:0] opcode,
	output[11:0] out

);
    
endmodule
